
interface dut_prm_if();
    bit             param_a, param_b, param_c;
endinterface

