
interface dut_out_if(input clk);
    logic           x, y, z;
endinterface

