
interface sig_if(input clk, rst_n);
    bit [0:2]   sig;
endinterface

