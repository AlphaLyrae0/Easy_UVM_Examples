
interface xyz_if(input clk, rst_n);
    logic           x, y, z;
endinterface

